module SPR(SR,Lo,Hi,clk);
  output [8:0] SR;
  output [15:0] Lo;
  output [15:0] Hi;
  input clk;
 
endmodule
